`timescale 1ns/1ps

module test_cbfp_tb;

    parameter array_size    = 16;
    parameter din_size      = 23;
    parameter dout_size     = 11;
    parameter buffer_depth  = 64;
    parameter array_num     = 4;
    parameter total_inputs  = 512;

    logic clk, rstn, valid_in;
    logic signed [din_size-1:0] din_re_p [0:array_size-1];
    logic signed [din_size-1:0] dout_re_p [0:array_size-1];
    logic [din_size-1:0] zero_cnt [0:array_num-1];

    integer file, r, i, j;
    integer data_array [0:total_inputs-1];
    string line;

    // DUT 연결
    test_cbfp #(
        .array_size(array_size),
        .din_size(din_size),
        .dout_size(dout_size),
        .buffer_depth(buffer_depth)
    ) uut (
        .clk(clk),
        .rstn(rstn),
        .valid_in(valid_in),
        .din_re_p(din_re_p),
        .dout_re_p(dout_re_p),
        .zero_cnt(zero_cnt)
    );

    // Clock generation (250MHz)
    always #2 clk = ~clk;

    initial begin
        $display("Start Simulation");

        clk = 0;
        rstn = 0;
        valid_in = 0;

        // 입력 초기화
        for (i = 0; i < array_size; i++) begin
            din_re_p[i] = 0;
        end

        // ===== 텍스트 파일 열기 =====
        file = $fopen("bfly02_tmp_fixed_real.txt", "r");
        if (file == 0) begin
            $display("Failed to open input file.");
            $finish;
        end

        // ===== 데이터 읽기 (최대 128개) =====
        for (i = 0; i < total_inputs; i++) begin
            r = $fscanf(file, "%d\n", data_array[i]);
        end
        $fclose(file);

        // ===== Reset =====
        #20;
        rstn = 1;
        #10;

        // ===== Phase 1: 첫 64개 입력 (4클럭 동안 16개씩) =====
        for (i = 192; i < 256; i += 16) begin
            valid_in = 1;
            for (j = 0; j < 16; j++) begin
                din_re_p[j] = data_array[i + j];
            end
            #4;
        end

        // ===== Phase 2: 입력 없음 (4클럭 동안 모두 0) =====
        for (i = 0; i < 4; i++) begin
            valid_in = 0;
            for (j = 0; j < 16; j++) begin
                din_re_p[j] = 0;
            end
            #4;
        end

        // ===== Phase 2: 다음 64개 입력 (4클럭 동안 16개씩) =====
        for (i = 256; i < 320; i += 16) begin
            valid_in = 1;
            for (j = 0; j < 16; j++) begin
                din_re_p[j] = data_array[i + j];
            end
            #4;
        end

        // ===== Phase 3: 입력 없음 (4클럭 동안 모두 0) =====
        for (i = 0; i < 4; i++) begin
            valid_in = 0;
            for (j = 0; j < 16; j++) begin
                din_re_p[j] = 0;
            end
            #4;
        end

        // ===== Phase 3: 다음 64개 입력 (4클럭 동안 16개씩) =====
        for (i = 320; i < 384; i += 16) begin
            valid_in = 1;
            for (j = 0; j < 16; j++) begin
                din_re_p[j] = data_array[i + j];
            end
            #4;
        end

        // ===== Phase 3: 입력 없음 (4클럭 동안 모두 0) =====
        for (i = 0; i < 4; i++) begin
            valid_in = 0;
            for (j = 0; j < 16; j++) begin
                din_re_p[j] = 0;
            end
            #4;
        end

        // ===== Phase 3: 다음 64개 입력 (4클럭 동안 16개씩) =====
        for (i = 384; i < 448; i += 16) begin
            valid_in = 1;
            for (j = 0; j < 16; j++) begin
                din_re_p[j] = data_array[i + j];
            end
            #4;
        end

        // 입력 종료
        valid_in = 0;

        // ===== 추가 시뮬레이션 시간 확보 =====
        #100;

        $display("Simulation End");
        $finish;
    end
endmodule
