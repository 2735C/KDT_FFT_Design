function automatic logic [4:0] count_min_lzc_23bit(input logic signed [22:0] din [0:15]);
    logic [4:0] lzc [0:15];
    logic [4:0] min_val = 21;

    for (int i = 0; i < 16; i++) begin
        lzc[i] =(din[i][21:0]  == 22'd0 && din[i][22] == 1'b0) ? 22 :
                (din[i][21:1]  == 21'd0 && din[i][22] == 1'b0) ? 21 :
                (din[i][21:2]  == 20'd0 && din[i][22] == 1'b0) ? 20 :
                (din[i][21:3]  == 19'd0 && din[i][22] == 1'b0) ? 19 :
                (din[i][21:4]  == 18'd0 && din[i][22] == 1'b0) ? 18 :
                (din[i][21:5]  == 17'd0 && din[i][22] == 1'b0) ? 17 :
                (din[i][21:6]  == 16'd0 && din[i][22] == 1'b0) ? 16 :
                (din[i][21:7]  == 15'd0 && din[i][22] == 1'b0) ? 15 :
                (din[i][21:8]  == 14'd0 && din[i][22] == 1'b0) ? 14 :
                (din[i][21:9]  == 13'd0 && din[i][22] == 1'b0) ? 13 :
                (din[i][21:10] == 12'd0 && din[i][22] == 1'b0) ? 12 :
                (din[i][21:11] == 11'd0 && din[i][22] == 1'b0) ? 11 :
                (din[i][21:12] == 10'd0 && din[i][22] == 1'b0) ? 10 :
                (din[i][21:13] == 9'd0  && din[i][22] == 1'b0) ? 9  :
                (din[i][21:14] == 8'd0  && din[i][22] == 1'b0) ? 8  :
                (din[i][21:15] == 7'd0  && din[i][22] == 1'b0) ? 7  :
                (din[i][21:16] == 6'd0  && din[i][22] == 1'b0) ? 6  :
                (din[i][21:17] == 5'd0  && din[i][22] == 1'b0) ? 5  :
                (din[i][21:18] == 4'd0  && din[i][22] == 1'b0) ? 4  :
                (din[i][21:19] == 3'd0  && din[i][22] == 1'b0) ? 3  :
                (din[i][21:20] == 2'd0  && din[i][22] == 1'b0) ? 2  :
                (din[i][21]    == 1'b0  && din[i][22] == 1'b0) ? 1  : 
                (din[i][21:0]  == 22'h3FFFFF && din[i][22] == 1'b1) ? 22 :
                (din[i][21:1]  == 21'h1FFFFF && din[i][22] == 1'b1) ? 21 :
                (din[i][21:2]  == 20'hFFFFF  && din[i][22] == 1'b1) ? 20 :
                (din[i][21:3]  == 19'h7FFFF  && din[i][22] == 1'b1) ? 19 :
                (din[i][21:4]  == 18'h3FFFF  && din[i][22] == 1'b1) ? 18 :
                (din[i][21:5]  == 17'h1FFFF  && din[i][22] == 1'b1) ? 17 :
                (din[i][21:6]  == 16'hFFFF   && din[i][22] == 1'b1) ? 16 :
                (din[i][21:7]  == 15'h7FFF   && din[i][22] == 1'b1) ? 15 :
                (din[i][21:8]  == 14'h3FFF   && din[i][22] == 1'b1) ? 14 :
                (din[i][21:9]  == 13'h1FFF   && din[i][22] == 1'b1) ? 13 :
                (din[i][21:10] == 12'hFFF    && din[i][22] == 1'b1) ? 12 :
                (din[i][21:11] == 11'h7FF    && din[i][22] == 1'b1) ? 11 :
                (din[i][21:12] == 10'h3FF    && din[i][22] == 1'b1) ? 10 :
                (din[i][21:13] ==  9'h1FF    && din[i][22] == 1'b1) ? 9  :
                (din[i][21:14] ==  8'hFF     && din[i][22] == 1'b1) ? 8  :
                (din[i][21:15] ==  7'h7F     && din[i][22] == 1'b1) ? 7  :
                (din[i][21:16] ==  6'h3F     && din[i][22] == 1'b1) ? 6  :
                (din[i][21:17] ==  5'h1F     && din[i][22] == 1'b1) ? 5  :
                (din[i][21:18] ==  4'hF      && din[i][22] == 1'b1) ? 4  :
                (din[i][21:19] ==  3'h7      && din[i][22] == 1'b1) ? 3  :
                (din[i][21:20] ==  2'h3      && din[i][22] == 1'b1) ? 2  :
                (din[i][21]    ==  1'b1      && din[i][22] == 1'b1) ? 1  : 0;

        if (lzc[i] < min_val)
            min_val = lzc[i];
    end

    return min_val;
endfunction
